module ALU (Out, In1, In2, COut, CIn, Op);
parameter op_size = 4;
input [31:0] In1, In2;
input [op_size-1:0] Op;
input CIn;
output [31:0] Out;
output Cout;





endmodule