`timescale 1 ns / 1 ps

module my_test_decoder;
    