module ALU (ac, mbr, Op, clk);
parameter op_size = 4;
input clk;
input [15:0] ac;
input [op_size-1:0] Op;
inout [15:0] mbr;





endmodule