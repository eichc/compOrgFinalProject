module MAR ();
    
endmodule